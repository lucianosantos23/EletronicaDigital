module teclado_para_xs3_tb;
    reg  [9:0] in;
    wire [3:0] out;

    teclado_para_xs3 dut (.in(in),.out(out));
    initial begin
        $monitor("in = %b, out (XS-3) = %b", in, out);
        in = 10'b0000000001; #10; // 0 -> 0011
        in = 10'b0000000010; #10; // 1 -> 0100
        in = 10'b0000000100; #10; // 2 -> 0101
        in = 10'b0000001000; #10; // 3 -> 0110
        in = 10'b0000010000; #10; // 4 -> 0111
        in = 10'b0000100000; #10; // 5 -> 1000
        in = 10'b0001000000; #10; // 6 -> 1001
        in = 10'b0010000000; #10; // 7 -> 1010
        in = 10'b0100000000; #10; // 8 -> 1011
        in = 10'b1000000000; #10; // 9 -> 1100
        $stop;
    end
endmodule
